module imem(
  input wire [31:0] a,
  output reg [31:0] rd
);
  reg [31:0] RAM[63:0] = '{
    32'h00500113, 32'h00C00193, 32'hFF718393, 32'h0023E233,
    32'h0041F2B3, 32'h004282B3, 32'h02728863, 32'h0041A233,
    32'h00020463, 32'h00000293, 32'h0023A233, 32'h005203B3,
    32'h402383B3, 32'h0471AA23, 32'h06002103, 32'h005104B3,
    32'h008001EF, 32'h00100113, 32'h00910133, 32'h0221A023,
    32'h00210063,
    // Add zeros to match the size of RAM
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
    32'h00000008, 32'h00000004, 32'h000000012    
  };

  // Perform word-aligned read
  assign rd = RAM[a[31:2]];

endmodule
